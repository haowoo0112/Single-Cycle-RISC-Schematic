// Verilog test fixture created from schematic C:\Users\USER\Desktop\Single-Cycle-RISC-Schematic\Single-Cycle-RISC-Schematic\D_flip_flop_16_bit.sch - Fri Sep 09 21:41:57 2022

`timescale 1ns / 1ps

module D_flip_flop_16_bit_D_flip_flop_16_bit_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   D_flip_flop_16_bit UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
